library verilog;
use verilog.vl_types.all;
entity WB_STAGE is
    port(
        ALU_result      : in     vl_logic_vector(31 downto 0);
        MEM_result      : in     vl_logic_vector(31 downto 0);
        MEM_R_en        : in     vl_logic;
        \out\           : out    vl_logic_vector(31 downto 0)
    );
end WB_STAGE;
