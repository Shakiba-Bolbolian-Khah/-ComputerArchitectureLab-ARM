`timescale 1ns/1ns
module INSTRUCTION_MEMORY(
  input[31:0] PC, output reg [31:0] Instruction
);
	wire [9:0] address;
  reg [31:0] memoryData[0:255];
	
	initial begin
		memoryData[0] = 32'b11100011101000000000000000010100;
    memoryData[1] = 32'b11100011101000000001101000000001;
    memoryData[2] = 32'b11100011101000000010000100000011;
    memoryData[3] = 32'b11100000100100100011000000000010;
    memoryData[4] = 32'b11100000101000000100000000000000;
    memoryData[5] = 32'b11100000010001000101000100000100;
    memoryData[6] = 32'b11100000110000000110000010100000;
    memoryData[7] = 32'b11100001100001010111000101000010;
    memoryData[8] = 32'b11100000000001111000000000000011;
    memoryData[9] = 32'b11100001111000001001000000000110;
    memoryData[10] = 32'b11100000001001001010000000000101;
    memoryData[11] = 32'b11100001010110000000000000000110;
    memoryData[12] = 32'b00010000100000010001000000000001;
    memoryData[13] = 32'b11100001000110010000000000001000;
    memoryData[14] = 32'b00000000100000100010000000000010;
    memoryData[15] = 32'b11100011101000000000101100000001;
    memoryData[16] = 32'b11100100100000000001000000000000;
    memoryData[17] = 32'b11100100100100001011000000000000;
    memoryData[18] = 32'b11100100100000000010000000000100;
    memoryData[19] = 32'b11100100100000000011000000001000;
    memoryData[20] = 32'b11100100100000000100000000001101;
    memoryData[21] = 32'b11100100100000000101000000010000;
    memoryData[22] = 32'b11100100100000000110000000010100;
    memoryData[23] = 32'b11100100100100001010000000000100;
    memoryData[24] = 32'b11100100100000000111000000011000;
    memoryData[25] = 32'b11100011101000000001000000000100;
    memoryData[26] = 32'b11100011101000000010000000000000;
    memoryData[27] = 32'b11100011101000000011000000000000;
    memoryData[28] = 32'b11100000100000000100000100000011;
    memoryData[29] = 32'b11100100100101000101000000000000;
    memoryData[30] = 32'b11100100100101000110000000000100;
    memoryData[31] = 32'b11100001010101010000000000000110;
    memoryData[32] = 32'b11000100100001000110000000000000;
    memoryData[33] = 32'b11000100100001000101000000000100;
    memoryData[34] = 32'b11100010100000110011000000000001;
    memoryData[35] = 32'b11100011010100110000000000000011;
    memoryData[36] = 32'b10111010111111111111111111110111;
    memoryData[37] = 32'b11100010100000100010000000000001;
    memoryData[38] = 32'b11100001010100100000000000000001;
    memoryData[39] = 32'b10111010111111111111111111110011;
    memoryData[40] = 32'b11100100100100000001000000000000;
    memoryData[41] = 32'b11100100100100000010000000000100;
    memoryData[42] = 32'b11100100100100000011000000001000;
    memoryData[43] = 32'b11100100100100000100000000001100;
    memoryData[44] = 32'b11100100100100000101000000010000;
    memoryData[45] = 32'b11100100100100000110000000010100;
    memoryData[46] = 32'b11101010111111111111111111111111;
  end

	assign address = (PC[9:0] >> 2);

  always@(PC)begin
		Instruction <= memoryData[address];
  end
endmodule